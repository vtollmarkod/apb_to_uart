package environment_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "my_environment.sv" 
	//`include "my_virtual_sequence.sv"
	//`include "my_virtual_sequencer.sv"

endpackage:environment_pkg