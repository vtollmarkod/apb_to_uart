interface uart_interface (input rst, input clk);
	logic rx;
	logic tx;
endinterface