interface uart_interface (input rst, input uart_clk);
	logic rx;
	logic tx;
endinterface