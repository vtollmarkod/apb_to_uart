class my_virtual_sequence extends uvm_sequence;
	`uvm_object_utils (my_virtual_seq)
    `uvm_declare_p_sequencer (my_virtual_sequencer)
  	
  function new(string name);
    super.new(name);
  endfunction
  
  
  // Zavristi nakon pakovanja u paket
  
  
  
  
endclass:my_virtual_sequence