	`include "apb_interface.sv"
package apb_pkg;
    import uvm_pkg::*;
    `include "apb_sequence_item.sv" 
    `include "apb_sequencer.sv"
    `include "apb_sequence.sv"
    `include "apb_driver.sv"
	`include "apb_monitor.sv"
	`include "apb_agent.sv"	
    `include "my_enviroment.sv"
    `include "apb_tests.sv"


endpackage: apb_pkg